class dti_scoreboard extends uvm_scoreboard;
  
endclass : dti_scoreboard