`include "uvm.sv"
`include "uvm_macros.svh"
import  uvm_pkg::*;

`include "mem_interface.sv"
`include "mem_seq_item.sv"
`include "mem_sequence.sv"
`include "mem_sequencer.sv"
`include "mem_driver.sv"
`include "mem_monitor.sv"
`include "mem_agent.sv"
`include "mem_scoreboard.sv"
`include "mem_env.sv"

`include "mem_base_test.sv"
`include "mem_wr_rd_test.sv"